library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bin_bcd is
    port(
        bin : in integer range 0 to 9999;   -- número en binario
        d0  : out std_logic_vector(3 downto 0); -- unidades
        d1  : out std_logic_vector(3 downto 0); -- decenas
        d2  : out std_logic_vector(3 downto 0); -- centenas
        d3  : out std_logic_vector(3 downto 0)  -- millares
    );
end bin_bcd;

architecture arch_bin_bcd of bin_bcd is
    signal value : integer range 0 to 9999;
begin
    process(bin)
        variable temp : integer range 0 to 9999;
        variable u, d, c, m : integer range 0 to 9;
    begin
        value <= bin;
        temp := bin;

        -- Cálculo de cada dígito (división sucesiva)
        m := temp / 1000;        -- millares
        temp := temp mod 1000;

        c := temp / 100;         -- centenas
        temp := temp mod 100;

        d := temp / 10;          -- decenas
        u := temp mod 10;        -- unidades

        -- Asignación a salidas en std_logic_vector
        d3 <= std_logic_vector(to_unsigned(m, 4));
        d2 <= std_logic_vector(to_unsigned(c, 4));
        d1 <= std_logic_vector(to_unsigned(d, 4));
        d0 <= std_logic_vector(to_unsigned(u, 4));
    end process;
end arch_bin_bcd;
